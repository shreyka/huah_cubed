`timescale 1ns / 1ps
`default_nettype none

/*

Given data from one block and an XY position,
render that block.

*/
module get_pixel_color(
    );
endmodule

`default_nettype wire