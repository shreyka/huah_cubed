`timescale 1ns / 1ps
`default_nettype none

module top_level(
  input wire clk_100mhz //clock @ 100 mhz
  );

  

endmodule




`default_nettype wire
