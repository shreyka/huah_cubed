`timescale 1ns / 1ps
`default_nettype none

/*

Given data from one block and an XY position,
render that block.

*/
module does_ray_block_intersect(
    );
endmodule

`default_nettype wire